module switch_level_modeling (
    input a,b,c;
    output d;
);
    
endmodule